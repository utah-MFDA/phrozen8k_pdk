
MACRO pump_40px_0
  CLASS CORE ;
  ORIGIN  0 0 ;
  FOREIGN pump_40px_0 0 0 ;
  SIZE 300 BY 115 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN in_fluid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 24.5 58.5 25.5 59.5 ;
    END
  END in_fluid
  PIN out_fluid
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 274.5 58.5 275.5 59.5 ;
    END
  END out_fluid
  PIN a_in_air
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 89.5 21.5 90.5 22.5 ;
    END
  END a_in_air
  PIN a_out_air
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 89.5 95.5 90.5 96.5 ;
    END
  END a_out_air
  PIN b_in_air
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 149.5 21.5 150.5 22.5 ;
    END
  END b_in_air
  PIN b_out_air
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 149.5 95.5 150.5 96.5 ;
    END
  END b_out_air
  PIN c_in_air
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 209.5 21.5 210.5 22.5 ;
    END
  END c_in_air
  PIN c_out_air
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 209.5 95.5 210.5 96.5 ;
    END
  END c_out_air
  OBS
    LAYER met1 ;
      RECT 25 22 275 96 ;
    LAYER met2 ;
      RECT 25 22 275 96 ;
    LAYER met3 ;
      RECT 25 22 275 96 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END pump_40px_0
