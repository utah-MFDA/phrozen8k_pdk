
MACRO valve_80px_1
  CLASS CORE ;
  ORIGIN  0 0 ;
  FOREIGN valve_80px_1 0 0 ;
  SIZE 190 BY 190 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN in_fluid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 29.5 91.5 30.5 92.5 ;
    END
  END in_fluid
  PIN out_fluid
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 158.5 91.5 159.5 92.5 ;
    END
  END out_fluid
  PIN in_air
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93 24.5 94 25.5 ;
    END
  END in_air
  PIN out_air
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93 159.5 94 160.5 ;
    END
  END out_air
  OBS
    LAYER met1 ;
      RECT 30 25 159 160 ;
    LAYER met2 ;
      RECT 30 25 159 160 ;
    LAYER met3 ;
      RECT 30 25 159 160 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END valve_80px_1
